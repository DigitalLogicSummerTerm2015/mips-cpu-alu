module shifter(
    output [31:0] dout,
    input [31:0] A,
    input [31:0] B,
    input [1:0] ctrl
);



endmodule
