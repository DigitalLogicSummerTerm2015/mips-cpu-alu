module comparer(
    output [31:0] dout,
    input Z,
    input V,
    input N,
    input [3:1] ctrl
);



endmodule
