module comparer(
    output [31:0] dout,
    input Z,  // Zero.
    input V,  // Overflow.
    input N,  // Negative.
    input [3:1] ctrl
);



endmodule
