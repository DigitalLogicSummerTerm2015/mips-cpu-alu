module adder(
    output Z,
    output V,
    output N,
    output [31:0] dout,
    input [31:0] A,
    input [31:0] B,
    input ctrl,

);



endmodule
